*** static buffer ***
*
* ngSPICE AND2X1 cell
*
* SPICE3 file originally created from AND2X1.ext by Magic - technology: scmos
*
*
* Author: Jan Belohoubek, 01/2020
* jan.belohoubek@fit.cvut.cz
*
* https://users.fit.cvut.cz/~belohja4/
*
*
* **************************************

.subckt AND2X1 A B O VSS VDD

X1000 Y A VDD VDD VSS LaserTrig SUBCKT_PMOS beamDistance = beamDistanceTop ch_w=2u ch_l=0.2u mos_ad=0.8p mos_pd=3.4u mos_as=0.8p mos_ps=3.4u
X1001 VDD B Y VDD VSS LaserTrig SUBCKT_PMOS beamDistance = beamDistanceTop ch_w=2u ch_l=0.2u mos_ad=0.7p mos_pd=3.4u mos_as=0.7p mos_ps=3.4u
X1002 O Y VDD VDD VSS LaserTrig SUBCKT_PMOS beamDistance = beamDistanceTop ch_w=2u ch_l=0.2u mos_ad=0.7p mos_pd=3.4u mos_as=0.7p mos_ps=3.4u

* mos_ad/mos_as partioning is correct, but because of small 1:2 transistor size partitioning, the photocurrent simmulation is not completely correct
X1003 MIDDLE A Y VSS psubIn LaserTrig   SUBCKT_NMOS beamDistance = beamDistanceBot ch_w=2u ch_l=0.2u mos_ad=1.1p mos_pd=4.6u mos_as=0.3p  mos_ps=0u commonDrain = 0 commonSource = 1
X1004 VSS B MIDDLE VSS psubIn LaserTrig SUBCKT_NMOS beamDistance = beamDistanceBot ch_w=2u ch_l=0.2u mos_ad=0.3p mos_pd=5.2u mos_as=0.75p mos_ps=3u commonDrain = 1 commonSource = 1
X1005 O Y VSS VSS psubIn LaserTrig      SUBCKT_NMOS beamDistance = beamDistanceBot ch_w=1u ch_l=0.2u mos_ad=0.5p mos_pd=3u   mos_as=0.25p mos_ps=2u commonDrain = 0 commonSource = 1

* common NMOS substarte virtual node
XpsubIn psubIn VSS PSUB_IN

C0 Y MIDDLE 0.00fF
C1 O VSS 0.19fF
C2 O Y 0.46fF
C3 Y VSS 0.10fF
C4 O VDD 0.38fF
C5 Y A 0.06fF
C6 Y VDD 0.82fF
C7 Y B 0.33fF
C8 A VDD 0.20fF
C9 A B 0.26fF
C10 VDD B 0.25fF
C11 VSS VSS 0.19fF
C12 O VSS 0.14fF
C13 Y VSS 0.38fF
C14 B VSS 0.19fF
C15 A VSS 0.25fF
C16 VDD VSS 1.73fF

.ends


