*** TEST 002 ***
*
* ngSPICE test for PLS experiments
*
* Current direction demonstration
*
* Author: Jan Belohoubek, 01/2019
* jan.belohoubek@fit.cvut.cz
*
* https://users.fit.cvut.cz/~belohja4/
*
*
* **************************************

.include ../models.lib


* **************************************
* --- Test Parameters ---
* **************************************

* **************************************
* --- Test ---
* **************************************

R1 VSS VDD 100

* **************************************
* --- Simulation Settings ---
* **************************************

.tran .1ns 100ns

* **************************************
* --- Simulation Control ---
* **************************************

.control
    run
    plot i(vvss) i(vvdd)

    echo PASSED
    
.endc

.end
